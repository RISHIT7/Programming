library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity my_module is
    port (
        clk : in std_logic;
        rst : in std_logic;
        sig
    );
end my_module;

architecture rtl of my_module is

begin

end architecture;